library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
entity s298_hot is
  port(
    clock:  in  std_logic;
    input:  in  std_logic_vector(2 downto 0);
    output: out std_logic_vector(5 downto 0)
  );
end s298_hot;
architecture behaviour of s298_hot is
  constant s00000000000000: std_logic_vector(217 downto 0) := "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000001100000: std_logic_vector(217 downto 0) := "01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000001100010: std_logic_vector(217 downto 0) := "00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000001100011: std_logic_vector(217 downto 0) := "00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000001100001: std_logic_vector(217 downto 0) := "00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000001100000: std_logic_vector(217 downto 0) := "00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000001100001: std_logic_vector(217 downto 0) := "00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000001100000: std_logic_vector(217 downto 0) := "00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000001100011: std_logic_vector(217 downto 0) := "00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000001100010: std_logic_vector(217 downto 0) := "00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001001100011: std_logic_vector(217 downto 0) := "00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001001100010: std_logic_vector(217 downto 0) := "00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001001100000: std_logic_vector(217 downto 0) := "00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001001100001: std_logic_vector(217 downto 0) := "00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100001100011: std_logic_vector(217 downto 0) := "00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100001100010: std_logic_vector(217 downto 0) := "00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100001100001: std_logic_vector(217 downto 0) := "00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100001100000: std_logic_vector(217 downto 0) := "00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101001100010: std_logic_vector(217 downto 0) := "00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101001100011: std_logic_vector(217 downto 0) := "00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101001100000: std_logic_vector(217 downto 0) := "00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101001100001: std_logic_vector(217 downto 0) := "00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01101001100010: std_logic_vector(217 downto 0) := "00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01101001100011: std_logic_vector(217 downto 0) := "00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01101001100001: std_logic_vector(217 downto 0) := "00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01101001100000: std_logic_vector(217 downto 0) := "00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00010001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00010001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00010001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00010001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000000011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01100001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01100001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01100001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01100001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11101000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00011001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10010001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11000100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10101100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10100100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00100100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s11001100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001010010001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001010010000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001010010011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00001010010010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000010010000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000000011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000000011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000000011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10000000011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s00101001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001000011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001000011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001000011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10001000011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001000011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001000011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001000011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01001000011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000000011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000000011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000000011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
  constant s01000000011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
  constant s10011001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
  constant s00000001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
  constant s00000001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000";
  constant s00000001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000";
  constant s10001001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000";
  constant s10001001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000";
  constant s10001001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000";
  constant s10001001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000";
  constant s10011010010000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000";
  constant s10011010010001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000";
  constant s10011010010010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000";
  constant s10011010010011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000";
  constant s00000010010011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000";
  constant s00000010010010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000";
  constant s00000010010001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000";
  constant s10010010010011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000";
  constant s10010010010010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000";
  constant s10010010010000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000";
  constant s10010010010001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000";
  constant s10011100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
  constant s10011100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000";
  constant s10011100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000";
  constant s10011100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
  constant s00000100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000";
  constant s00000100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000";
  constant s00000100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000";
  constant s00000100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000";
  constant s11100001100001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
  constant s11100001100000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000";
  constant s11100001100010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000";
  constant s11100001100011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
  constant s10010000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000";
  constant s10010000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000";
  constant s10010000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000";
  constant s10010000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
  constant s00010000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000";
  constant s00010000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000";
  constant s00010000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000";
  constant s00010000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000";
  constant s11100000100111: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000";
  constant s11100000100110: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000";
  constant s11100000100100: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000";
  constant s11100000100101: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000";
  constant s01100100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000";
  constant s01100100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000";
  constant s01100100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000";
  constant s01100100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000";
  constant s11100100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000";
  constant s11100100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000";
  constant s11100100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000";
  constant s11100100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000";
  constant s00011100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000";
  constant s00011100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000";
  constant s00011100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000";
  constant s00011100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000";
  constant s00010100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000";
  constant s00010100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000";
  constant s00010100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000";
  constant s00010100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000";
  constant s11101100011001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000";
  constant s11101100011000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000";
  constant s11101100011010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000";
  constant s11101100011011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000";
  constant s01101100000000: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000";
  constant s01101100000001: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100";
  constant s01101100000011: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
  constant s01101100000010: std_logic_vector(217 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
  signal current_state, next_state: std_logic_vector(217 downto 0);
begin
  process(clock) begin
    if rising_edge(clock) then current_state <= next_state;
    end if;
  end process;
  process(input, current_state) begin
    next_state <= "--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------"; output <= "------";
    case current_state is
      when s00000000000000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10000001100010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10000001100011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10000001100001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10000001100000; output <= "000000";
        end if;
      when s00000001100000 =>
        if std_match(input, "000") then next_state <= s10000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10000001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10000001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10000001100011; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10000001100000 =>
        if std_match(input, "010") then next_state <= s01000001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01000001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01000001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01000001100001 =>
        if std_match(input, "001") then next_state <= s11001001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11001001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11001001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11001001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s11001001100011 =>
        if std_match(input, "000") then next_state <= s00100001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00100001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00100001100001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00100001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00100001100011 =>
        if std_match(input, "010") then next_state <= s10101001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10101001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10101001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10101001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10101001100010 =>
        if std_match(input, "000") then next_state <= s01101001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01101001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01101001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01101001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01101001100010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11101001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11101001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11101001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11101001100001; output <= "100001";
        end if;
      when s11101001100011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00010001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00010001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00010001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00010001100001; output <= "100001";
        end if;
      when s00010001100010 =>
        if std_match(input, "000") then next_state <= s10010100011010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10010100011011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10010100011000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10010100011001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "100001";
        end if;
      when s10010100011010 =>
        if std_match(input, "011") then next_state <= s00001100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00001100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00001100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00001100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s00001100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10000100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10000100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10000100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10000100011011; output <= "000000";
        end if;
      when s00000000011000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s10000001100010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s10000001100011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s10000001100000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s10000001100001; output <= "010100";
        end if;
      when s10000001100010 =>
        if std_match(input, "010") then next_state <= s01000001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01000001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01000001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01000001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01000001100011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11001001100001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11001001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11001001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11001001100010; output <= "100001";
        end if;
      when s11001001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00100001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00100001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00100001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00100001100010; output <= "100001";
        end if;
      when s00100001100000 =>
        if std_match(input, "001") then next_state <= s10100001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10100001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10100001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10100001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10100001100010 =>
        if std_match(input, "011") then next_state <= s01100001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01100001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01100001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01100001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01100001100001 =>
        if std_match(input, "011") then next_state <= s11101000100110; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11101000100111; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11101000100101; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11101000100100; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        end if;
      when s11101000100110 =>
        if std_match(input, "000") then next_state <= s00011000100110; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00011000100111; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00011000100101; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00011000100100; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s00011000100110 =>
        if std_match(input, "001") then next_state <= s10011000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10011000100101; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10011000100111; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10011000100110; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s10011000100100 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00000000100111; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00000000100110; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00000000100101; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s00000000100100 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10000001100010; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10000001100011; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10000001100000; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10000001100001; output <= "100010";
        end if;
      when s10000001100011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01001001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01001001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01001001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01001001100001; output <= "100001";
        end if;
      when s01001001100011 =>
        if std_match(input, "011") then next_state <= s11000001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11000001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11000001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11000001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s11000001100000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00100001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00100001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00100001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00100001100000; output <= "100001";
        end if;
      when s00100001100010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10100001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10100001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10100001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10100001100001; output <= "100001";
        end if;
      when s10100001100011 =>
        if std_match(input, "011") then next_state <= s01101001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01101001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01101001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01101001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01101001100000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11101001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11101001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11101001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11101001100000; output <= "100001";
        end if;
      when s11101001100010 =>
        if std_match(input, "011") then next_state <= s00011001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00011001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00011001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00011001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00011001100001 =>
        if std_match(input, "011") then next_state <= s10010001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10010001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10010001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10010001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10010001100010 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00001100000010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00001100000011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00001100000001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00001100000000; output <= "100001";
        end if;
      when s00001100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10001100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10001100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10001100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10001100011010; output <= "000000";
        end if;
      when s10001100011000 =>
        if std_match(input, "010") then next_state <= s01001100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s01001100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11000100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11000100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11000100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11000100011011; output <= "000000";
        end if;
      when s11000100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00101100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00101100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00101100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00101100000011; output <= "010100";
        end if;
      when s00101100000000 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10101100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10101100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10101100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10101100011011; output <= "000000";
        end if;
      when s00101100000001 =>
        if std_match(input, "001") then next_state <= s10100100011011; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10100100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10100100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10100100011000; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s00101100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10101100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10101100011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10101100011010; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10101100011011; output <= "000000";
        end if;
      when s00101100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10100100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10100100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10100100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10100100011010; output <= "000000";
        end if;
      when s11000100011000 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00100100000011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00100100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00100100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00100100000000; output <= "010100";
        end if;
      when s00100100000011 =>
        if std_match(input, "011") then next_state <= s10101100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10101100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10101100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10101100011011; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s00100100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10100100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10100100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10100100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10100100011010; output <= "000000";
        end if;
      when s00100100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10101100011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10101100011001; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10101100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10101100011011; output <= "000000";
        end if;
      when s00100100000000 =>
        if std_match(input, "000") then next_state <= s10100100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10100100011001; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10100100011011; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10100100011010; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s11000100011010 =>
        if std_match(input, "011") then next_state <= s00100100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00100100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00100100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00100100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s11000100011011 =>
        if std_match(input, "010") then next_state <= s00101100000010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00101100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00101100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00101100000001; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s01001100000000 =>
        if std_match(input, "000") then next_state <= s11001100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11001100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11001100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11001100011011; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s11001100011000 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00101100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00101100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00101100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00101100000011; output <= "010100";
        end if;
      when s11001100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00100100000001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00100100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00100100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00100100000010; output <= "010100";
        end if;
      when s11001100011010 =>
        if std_match(input, "000") then next_state <= s00101100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00101100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00101100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00101100000000; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s11001100011011 =>
        if std_match(input, "001") then next_state <= s00100100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00100100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00100100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00100100000010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s01001100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11001100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11001100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11001100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11001100011001; output <= "000000";
        end if;
      when s01001100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11000100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11000100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11000100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11000100011010; output <= "000000";
        end if;
      when s10001100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01000100000011; output <= "010100";
        end if;
      when s01000100000000 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11000100011011; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11000100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11000100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11000100011001; output <= "000000";
        end if;
      when s01000100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11001100011011; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11001100011010; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11001100011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11001100011001; output <= "000000";
        end if;
      when s01000100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11000100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11000100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11000100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11000100011010; output <= "000000";
        end if;
      when s01000100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11001100011001; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11001100011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11001100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11001100011010; output <= "000000";
        end if;
      when s10001100011011 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000100000010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000100000011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01000100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000100000000; output <= "010100";
        end if;
      when s10001100011010 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01001100000011; output <= "010100";
        end if;
      when s00001100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10000100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10000100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10000100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10000100011011; output <= "000000";
        end if;
      when s10000100011000 =>
        if std_match(input, "001") then next_state <= s01000100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000100000011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000100000001; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s10000100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001100000011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001100000001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01001100000000; output <= "010100";
        end if;
      when s10000100011010 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01000100000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000100000011; output <= "010100";
        end if;
      when s10000100011011 =>
        if std_match(input, "011") then next_state <= s01001100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001100000001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01001100000010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s00001100000000 =>
        if std_match(input, "011") then next_state <= s10001100011011; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10001100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10001100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10001100011001; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s10010001100011 =>
        if std_match(input, "001") then next_state <= s00001100000001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00001100000000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00001100000010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00001100000011; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "100001";
        end if;
      when s10010001100001 =>
        if std_match(input, "000") then next_state <= s00001010010001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00001010010000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00001010010011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00001010010010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000010010000; output <= "100001";
        end if;
      when s00001010010001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s10000000011010; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10000000011011; output <= "001100";
        elsif std_match(input, "000") then next_state <= s10000000011001; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10000000011000; output <= "001100";
        end if;
      when s10000000011010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000001100010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000001100011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01000001100000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000001100001; output <= "010100";
        end if;
      when s01000001100010 =>
        if std_match(input, "000") then next_state <= s11000001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11000001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11000001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11000001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s11000001100010 =>
        if std_match(input, "000") then next_state <= s00100001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00100001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00100001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00100001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00100001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10101001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10101001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10101001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10101001100000; output <= "100001";
        end if;
      when s11000001100011 =>
        if std_match(input, "010") then next_state <= s00101001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00101001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00101001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00101001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00101001100010 =>
        if std_match(input, "001") then next_state <= s10101001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10101001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10101001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10101001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00101001100011 =>
        if std_match(input, "011") then next_state <= s10100001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10100001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10100001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10100001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00101001100000 =>
        if std_match(input, "001") then next_state <= s10101001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10101001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10101001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10101001100000; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00101001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10100001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10100001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10100001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10100001100001; output <= "100001";
        end if;
      when s11000001100001 =>
        if std_match(input, "001") then next_state <= s00101001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00101001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00101001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00101001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01000001100000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11000001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11000001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11000001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11000001100011; output <= "100001";
        end if;
      when s10000000011011 =>
        if std_match(input, "001") then next_state <= s01001001100001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001001100000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01001001100010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001001100011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        end if;
      when s01001001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11000001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11000001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11000001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11000001100010; output <= "100001";
        end if;
      when s01001001100000 =>
        if std_match(input, "010") then next_state <= s11001001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11001001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11001001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11001001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s11001001100000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00101001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00101001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00101001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00101001100001; output <= "100001";
        end if;
      when s11001001100010 =>
        if std_match(input, "001") then next_state <= s00101001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00101001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00101001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00101001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01001001100010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11001001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11001001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11001001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11001001100011; output <= "100001";
        end if;
      when s10000000011001 =>
        if std_match(input, "010") then next_state <= s01001001100000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001001100001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001001100011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001001100010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        end if;
      when s10000000011000 =>
        if std_match(input, "000") then next_state <= s01000001100000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000001100001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000001100011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01000001100010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        end if;
      when s00001010010000 =>
        if std_match(input, "000") then next_state <= s10001000011000; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10001000011001; output <= "001100";
        elsif std_match(input, "011") then next_state <= s10001000011011; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10001000011010; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "001100";
        end if;
      when s10001000011000 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001000011011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001000011010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01001000011001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01001000011000; output <= "010100";
        end if;
      when s01001000011011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11000001100011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11000001100010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11000001100001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11000001100000; output <= "010100";
        end if;
      when s01001000011010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11001001100010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11001001100011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11001001100000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11001001100001; output <= "010100";
        end if;
      when s01001000011001 =>
        if std_match(input, "001") then next_state <= s11000001100011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11000001100010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11000001100001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11000001100000; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        end if;
      when s01001000011000 =>
        if std_match(input, "010") then next_state <= s11001001100001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11001001100000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11001001100011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11001001100010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        end if;
      when s10001000011001 =>
        if std_match(input, "001") then next_state <= s01000000011011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000000011010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000000011001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000000011000; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "010100";
        end if;
      when s01000000011011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11001001100001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11001001100000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11001001100010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11001001100011; output <= "010100";
        end if;
      when s01000000011010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11000001100011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11000001100010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11000001100000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11000001100001; output <= "010100";
        end if;
      when s01000000011001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11001001100011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11001001100010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11001001100001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11001001100000; output <= "010100";
        end if;
      when s01000000011000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s11000001100000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s11000001100001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s11000001100010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s11000001100011; output <= "010100";
        end if;
      when s10001000011011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01000000011010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01000000011011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01000000011001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01000000011000; output <= "010100";
        end if;
      when s10001000011010 =>
        if std_match(input, "000") then next_state <= s01001000011010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01001000011011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01001000011001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01001000011000; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "010100";
        end if;
      when s00001010010011 =>
        if std_match(input, "010") then next_state <= s10000000011010; output <= "001100";
        elsif std_match(input, "000") then next_state <= s10000000011011; output <= "001100";
        elsif std_match(input, "011") then next_state <= s10000000011000; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10000000011001; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "001100";
        end if;
      when s00001010010010 =>
        if std_match(input, "000") then next_state <= s10001000011010; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10001000011011; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10001000011000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s10001000011001; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "001100";
        end if;
      when s00000010010000 =>
        if std_match(input, "011") then next_state <= s10000001100011; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10000001100010; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10000001100001; output <= "001100";
        elsif std_match(input, "000") then next_state <= s10000001100000; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "001100";
        end if;
      when s10000001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01001001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01001001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01001001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01001001100000; output <= "100001";
        end if;
      when s10010001100000 =>
        if std_match(input, "010") then next_state <= s00001010010001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00001010010000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00001010010011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00001010010010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000010010000; output <= "100001";
        end if;
      when s00011001100000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10011001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10011001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10011001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10011001100010; output <= "100001";
        end if;
      when s10011001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00000001100001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00000001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00000001100011; output <= "100001";
        end if;
      when s00000001100001 =>
        if std_match(input, "010") then next_state <= s10001001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10001001100001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10001001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10001001100011; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10001001100000 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01001000011010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01001000011011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01001000011001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01001000011000; output <= "100001";
        end if;
      when s10001001100001 =>
        if std_match(input, "000") then next_state <= s01000000011001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01000000011000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01000000011010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01000000011011; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "100001";
        end if;
      when s10001001100010 =>
        if std_match(input, "010") then next_state <= s01001000011011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01001000011010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01001000011000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01001000011001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "100001";
        end if;
      when s10001001100011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01000000011011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01000000011010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01000000011000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01000000011001; output <= "100001";
        end if;
      when s00000001100010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10000001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10000001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10000001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10000001100000; output <= "100001";
        end if;
      when s00000001100011 =>
        if std_match(input, "011") then next_state <= s10001001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10001001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10001001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10001001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10011001100000 =>
        if std_match(input, "1-1") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00000001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00000001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00000001100001; output <= "100001";
        elsif std_match(input, "110") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "-00") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10011001100011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00000001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00000001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00000001100001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10011001100010 =>
        if std_match(input, "000") then next_state <= s00000001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00000001100011; output <= "100001";
        elsif std_match(input, "1-0") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "1-1") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00000001100001; output <= "100001";
        end if;
      when s00011001100011 =>
        if std_match(input, "011") then next_state <= s10010001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10010001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10010001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10010001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00011001100010 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10011001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10011001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10011001100010; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10011001100011; output <= "100001";
        end if;
      when s11101001100001 =>
        if std_match(input, "000") then next_state <= s00010001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00010001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00010001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00010001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s00010001100001 =>
        if std_match(input, "1--") then next_state <= s00000010010000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10011010010000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10011010010001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10011010010010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10011010010011; output <= "100001";
        end if;
      when s10011010010000 =>
        if std_match(input, "011") then next_state <= s00000010010011; output <= "001100";
        elsif std_match(input, "001") then next_state <= s00000010010010; output <= "001100";
        elsif std_match(input, "1-1") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "1-0") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "010") then next_state <= s00000010010001; output <= "001100";
        elsif std_match(input, "000") then next_state <= s00000010010000; output <= "001100";
        end if;
      when s00000010010011 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s10001001100000; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10001001100001; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10001001100010; output <= "001100";
        elsif std_match(input, "000") then next_state <= s10001001100011; output <= "001100";
        end if;
      when s00000010010010 =>
        if std_match(input, "011") then next_state <= s10000001100001; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10000001100000; output <= "001100";
        elsif std_match(input, "000") then next_state <= s10000001100010; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10000001100011; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "001100";
        end if;
      when s00000010010001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "001100";
        elsif std_match(input, "000") then next_state <= s10001001100001; output <= "001100";
        elsif std_match(input, "010") then next_state <= s10001001100000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s10001001100010; output <= "001100";
        elsif std_match(input, "001") then next_state <= s10001001100011; output <= "001100";
        end if;
      when s10011010010001 =>
        if std_match(input, "001") then next_state <= s00000010010011; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00000010010010; output <= "001100";
        elsif std_match(input, "1-1") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "000") then next_state <= s00000010010001; output <= "001100";
        elsif std_match(input, "100") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "-10") then next_state <= s00000010010000; output <= "001100";
        end if;
      when s10011010010010 =>
        if std_match(input, "000") then next_state <= s00000010010010; output <= "001100";
        elsif std_match(input, "010") then next_state <= s00000010010011; output <= "001100";
        elsif std_match(input, "1-0") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "111") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00000010010001; output <= "001100";
        elsif std_match(input, "-01") then next_state <= s00000010010000; output <= "001100";
        end if;
      when s10011010010011 =>
        if std_match(input, "1--") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00000010010000; output <= "001100";
        elsif std_match(input, "001") then next_state <= s00000010010001; output <= "001100";
        elsif std_match(input, "000") then next_state <= s00000010010011; output <= "001100";
        elsif std_match(input, "010") then next_state <= s00000010010010; output <= "001100";
        end if;
      when s00010001100000 =>
        if std_match(input, "011") then next_state <= s10010010010011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10010010010010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10010010010000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10010010010001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000010010000; output <= "100001";
        end if;
      when s10010010010011 =>
        if std_match(input, "000") then next_state <= s00001100000011; output <= "001100";
        elsif std_match(input, "010") then next_state <= s00001100000010; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00001100000000; output <= "001100";
        elsif std_match(input, "001") then next_state <= s00001100000001; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "001100";
        end if;
      when s10010010010010 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "001100";
        elsif std_match(input, "001") then next_state <= s00001100000000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00001100000001; output <= "001100";
        elsif std_match(input, "000") then next_state <= s00001100000010; output <= "001100";
        elsif std_match(input, "010") then next_state <= s00001100000011; output <= "001100";
        end if;
      when s10010010010000 =>
        if std_match(input, "010") then next_state <= s00001010010001; output <= "001100";
        elsif std_match(input, "000") then next_state <= s00001010010000; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00001010010011; output <= "001100";
        elsif std_match(input, "001") then next_state <= s00001010010010; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000010010000; output <= "001100";
        end if;
      when s10010010010001 =>
        if std_match(input, "010") then next_state <= s00001010010000; output <= "001100";
        elsif std_match(input, "000") then next_state <= s00001010010001; output <= "001100";
        elsif std_match(input, "011") then next_state <= s00001010010010; output <= "001100";
        elsif std_match(input, "001") then next_state <= s00001010010011; output <= "001100";
        elsif std_match(input, "1--") then next_state <= s00000010010000; output <= "001100";
        end if;
      when s00010001100011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s10011100011000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s10011100011001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s10011100011011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s10011100011010; output <= "100001";
        end if;
      when s10011100011000 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00000100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00000100000011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00000100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00000100000001; output <= "010100";
        end if;
      when s00000100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10000100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10000100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10000100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10000100011000; output <= "000000";
        end if;
      when s00000100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10001100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10001100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10001100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10001100011010; output <= "000000";
        end if;
      when s00000100000000 =>
        if std_match(input, "001") then next_state <= s10000100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10000100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10000100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10000100011001; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s00000100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10001100011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10001100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10001100011011; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10001100011010; output <= "000000";
        end if;
      when s10011100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00000100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00000100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00000100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00000100000001; output <= "010100";
        end if;
      when s10011100011011 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00000100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00000100000001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00000100000010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00000100000011; output <= "010100";
        end if;
      when s10011100011010 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00000100000011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00000100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00000100000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00000100000001; output <= "010100";
        end if;
      when s11101001100000 =>
        if std_match(input, "011") then next_state <= s00011001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00011001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00011001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00011001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01101001100001 =>
        if std_match(input, "000") then next_state <= s11100001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11100001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11100001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11100001100011; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s11100001100001 =>
        if std_match(input, "001") then next_state <= s00011000100111; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00011000100110; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00011000100100; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00011000100101; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        end if;
      when s00011000100111 =>
        if std_match(input, "000") then next_state <= s10010000100111; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10010000100110; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10010000100101; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10010000100100; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s10010000100111 =>
        if std_match(input, "000") then next_state <= s00001100000011; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00001100000010; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00001100000001; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00001100000000; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "100010";
        end if;
      when s10010000100110 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00001100000010; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00001100000011; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00001100000000; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00001100000001; output <= "100010";
        end if;
      when s10010000100101 =>
        if std_match(input, "010") then next_state <= s00001010010000; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00001010010001; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00001010010011; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00001010010010; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000010010000; output <= "100010";
        end if;
      when s10010000100100 =>
        if std_match(input, "1--") then next_state <= s00000010010000; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00001010010000; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00001010010001; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00001010010011; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00001010010010; output <= "100010";
        end if;
      when s00011000100100 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10011000100110; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10011000100111; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10011000100101; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10011000100100; output <= "100010";
        end if;
      when s10011000100110 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00000000100101; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00000000100110; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00000000100111; output <= "100010";
        end if;
      when s00000000100101 =>
        if std_match(input, "001") then next_state <= s10001001100011; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10001001100010; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10001001100000; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10001001100001; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100010";
        end if;
      when s00000000100110 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10000001100011; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10000001100010; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10000001100001; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10000001100000; output <= "100010";
        end if;
      when s00000000100111 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10001001100001; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10001001100000; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10001001100010; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10001001100011; output <= "100010";
        end if;
      when s10011000100111 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00000000100111; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00000000100110; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00000000100101; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s10011000100101 =>
        if std_match(input, "011") then next_state <= s00000000100110; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00000000100111; output <= "100010";
        elsif std_match(input, "1-1") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "1-0") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00000000100101; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s00011000100101 =>
        if std_match(input, "000") then next_state <= s10010000100101; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10010000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10010000100110; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10010000100111; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s11100001100000 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00010000100100; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00010000100101; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00010000100110; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00010000100111; output <= "100001";
        end if;
      when s00010000100100 =>
        if std_match(input, "1--") then next_state <= s00000010010000; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10010010010010; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10010010010011; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10010010010000; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10010010010001; output <= "100010";
        end if;
      when s00010000100101 =>
        if std_match(input, "1--") then next_state <= s00000010010000; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10011010010000; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10011010010001; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10011010010011; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10011010010010; output <= "100010";
        end if;
      when s00010000100110 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10010100011000; output <= "100010";
        elsif std_match(input, "011") then next_state <= s10010100011001; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10010100011011; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10010100011010; output <= "100010";
        end if;
      when s10010100011000 =>
        if std_match(input, "010") then next_state <= s00001100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00001100000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00001100000011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00001100000010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s10010100011001 =>
        if std_match(input, "010") then next_state <= s00001100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00001100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00001100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00001100000010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s10010100011011 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00001100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00001100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00001100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00001100000001; output <= "010100";
        end if;
      when s00010000100111 =>
        if std_match(input, "011") then next_state <= s10011100011000; output <= "100010";
        elsif std_match(input, "001") then next_state <= s10011100011001; output <= "100010";
        elsif std_match(input, "010") then next_state <= s10011100011010; output <= "100010";
        elsif std_match(input, "000") then next_state <= s10011100011011; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "100010";
        end if;
      when s11100001100010 =>
        if std_match(input, "001") then next_state <= s00010000100100; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00010000100101; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00010000100111; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00010000100110; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        end if;
      when s11100001100011 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        elsif std_match(input, "001") then next_state <= s00011000100101; output <= "100001";
        elsif std_match(input, "011") then next_state <= s00011000100100; output <= "100001";
        elsif std_match(input, "000") then next_state <= s00011000100111; output <= "100001";
        elsif std_match(input, "010") then next_state <= s00011000100110; output <= "100001";
        end if;
      when s01101001100011 =>
        if std_match(input, "000") then next_state <= s11100001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11100001100010; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11100001100000; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11100001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10100001100000 =>
        if std_match(input, "011") then next_state <= s01100001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01100001100010; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01100001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01100001100001; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s01100001100011 =>
        if std_match(input, "010") then next_state <= s11101000100110; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11101000100111; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11101000100100; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11101000100101; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        end if;
      when s11101000100111 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00010000100110; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00010000100111; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00010000100101; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00010000100100; output <= "100010";
        end if;
      when s11101000100100 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00011000100100; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00011000100101; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00011000100111; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00011000100110; output <= "100010";
        end if;
      when s11101000100101 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00010000100110; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00010000100111; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00010000100101; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00010000100100; output <= "100010";
        end if;
      when s01100001100010 =>
        if std_match(input, "010") then next_state <= s11100000100111; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11100000100110; output <= "100001";
        elsif std_match(input, "001") then next_state <= s11100000100100; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11100000100101; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        end if;
      when s11100000100111 =>
        if std_match(input, "011") then next_state <= s00011000100100; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00011000100101; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00011000100110; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00011000100111; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s11100000100110 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00010000100110; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00010000100111; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00010000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00010000100101; output <= "100010";
        end if;
      when s11100000100100 =>
        if std_match(input, "011") then next_state <= s00010000100111; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00010000100110; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00010000100100; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00010000100101; output <= "100010";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        end if;
      when s11100000100101 =>
        if std_match(input, "1--") then next_state <= s00000000100100; output <= "100010";
        elsif std_match(input, "011") then next_state <= s00011000100110; output <= "100010";
        elsif std_match(input, "001") then next_state <= s00011000100111; output <= "100010";
        elsif std_match(input, "000") then next_state <= s00011000100101; output <= "100010";
        elsif std_match(input, "010") then next_state <= s00011000100100; output <= "100010";
        end if;
      when s01100001100000 =>
        if std_match(input, "001") then next_state <= s11100000100110; output <= "100001";
        elsif std_match(input, "011") then next_state <= s11100000100111; output <= "100001";
        elsif std_match(input, "000") then next_state <= s11100000100100; output <= "100001";
        elsif std_match(input, "010") then next_state <= s11100000100101; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000000100100; output <= "100001";
        end if;
      when s10100001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01101001100010; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01101001100011; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01101001100001; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01101001100000; output <= "100001";
        end if;
      when s10101001100011 =>
        if std_match(input, "001") then next_state <= s01100001100001; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01100001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01100001100011; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01100001100010; output <= "100001";
        elsif std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        end if;
      when s10101001100000 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01101001100001; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01101001100000; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01101001100011; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01101001100010; output <= "100001";
        end if;
      when s10101001100001 =>
        if std_match(input, "1--") then next_state <= s00000001100000; output <= "100001";
        elsif std_match(input, "010") then next_state <= s01100001100000; output <= "100001";
        elsif std_match(input, "000") then next_state <= s01100001100001; output <= "100001";
        elsif std_match(input, "001") then next_state <= s01100001100011; output <= "100001";
        elsif std_match(input, "011") then next_state <= s01100001100010; output <= "100001";
        end if;
      when s10100100011000 =>
        if std_match(input, "001") then next_state <= s01100100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01100100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01100100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01100100000000; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s01100100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11100100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11100100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11100100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11100100011000; output <= "000000";
        end if;
      when s11100100011011 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00011100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00011100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00011100000010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00011100000011; output <= "010100";
        end if;
      when s00011100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10010100011011; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10010100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10010100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10010100011000; output <= "000000";
        end if;
      when s00011100000000 =>
        if std_match(input, "000") then next_state <= s10011100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10011100011001; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10011100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10011100011011; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s00011100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10011100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10011100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10011100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10011100011001; output <= "000000";
        end if;
      when s00011100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10010100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10010100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10010100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10010100011010; output <= "000000";
        end if;
      when s11100100011010 =>
        if std_match(input, "001") then next_state <= s00010100000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00010100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00010100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00010100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s00010100000000 =>
        if std_match(input, "010") then next_state <= s10010100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10010100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10010100011011; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10010100011010; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s00010100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10011100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10011100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10011100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10011100011000; output <= "000000";
        end if;
      when s00010100000010 =>
        if std_match(input, "001") then next_state <= s10010100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10010100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s10010100011010; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10010100011011; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s00010100000011 =>
        if std_match(input, "000") then next_state <= s10011100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s10011100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s10011100011001; output <= "000000";
        elsif std_match(input, "011") then next_state <= s10011100011000; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s11100100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00011100000001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00011100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00011100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00011100000010; output <= "010100";
        end if;
      when s11100100011000 =>
        if std_match(input, "010") then next_state <= s00010100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00010100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00010100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00010100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s01100100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11101100011001; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11101100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11101100011010; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11101100011011; output <= "000000";
        end if;
      when s11101100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00010100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00010100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00010100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00010100000001; output <= "010100";
        end if;
      when s11101100011000 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00011100000010; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00011100000011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00011100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00011100000001; output <= "010100";
        end if;
      when s11101100011010 =>
        if std_match(input, "011") then next_state <= s00011100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00011100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00011100000011; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00011100000010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s11101100011011 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s00010100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s00010100000010; output <= "010100";
        elsif std_match(input, "001") then next_state <= s00010100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s00010100000000; output <= "010100";
        end if;
      when s01100100000001 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11101100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11101100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11101100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11101100011011; output <= "000000";
        end if;
      when s01100100000000 =>
        if std_match(input, "000") then next_state <= s11100100011000; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11100100011001; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11100100011011; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11100100011010; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s10100100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01101100000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01101100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01101100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01101100000010; output <= "010100";
        end if;
      when s01101100000000 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11101100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11101100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11101100011001; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11101100011000; output <= "000000";
        end if;
      when s01101100000001 =>
        if std_match(input, "011") then next_state <= s11100100011010; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11100100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11100100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11100100011000; output <= "000000";
        elsif std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        end if;
      when s01101100000011 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11100100011011; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11100100011010; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11100100011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11100100011001; output <= "000000";
        end if;
      when s01101100000010 =>
        if std_match(input, "1--") then next_state <= s00000000011000; output <= "000000";
        elsif std_match(input, "001") then next_state <= s11101100011000; output <= "000000";
        elsif std_match(input, "011") then next_state <= s11101100011001; output <= "000000";
        elsif std_match(input, "010") then next_state <= s11101100011011; output <= "000000";
        elsif std_match(input, "000") then next_state <= s11101100011010; output <= "000000";
        end if;
      when s10100100011011 =>
        if std_match(input, "011") then next_state <= s01101100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01101100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01101100000011; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01101100000010; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s10100100011010 =>
        if std_match(input, "001") then next_state <= s01100100000000; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01100100000001; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01100100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01100100000011; output <= "010100";
        elsif std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        end if;
      when s10101100011000 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01101100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01101100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01101100000011; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01101100000010; output <= "010100";
        end if;
      when s10101100011001 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01100100000001; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01100100000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01100100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01100100000010; output <= "010100";
        end if;
      when s10101100011010 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01101100000010; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01101100000011; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01101100000001; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01101100000000; output <= "010100";
        end if;
      when s10101100011011 =>
        if std_match(input, "1--") then next_state <= s00000000000000; output <= "010100";
        elsif std_match(input, "001") then next_state <= s01100100000001; output <= "010100";
        elsif std_match(input, "011") then next_state <= s01100100000000; output <= "010100";
        elsif std_match(input, "010") then next_state <= s01100100000010; output <= "010100";
        elsif std_match(input, "000") then next_state <= s01100100000011; output <= "010100";
        end if;
      when others => next_state <= "--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------"; output <= "------";
    end case;
  end process;
end behaviour;
