library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
entity tbk_rnd is
  port(
    clock:  in  std_logic;
    input:  in  std_logic_vector(5 downto 0);
    output: out std_logic_vector(2 downto 0)
  );
end tbk_rnd;
architecture behaviour of tbk_rnd is
  constant st0: std_logic_vector(4 downto 0) := "11101";
  constant st16: std_logic_vector(4 downto 0) := "00010";
  constant st1: std_logic_vector(4 downto 0) := "11011";
  constant st2: std_logic_vector(4 downto 0) := "11110";
  constant st3: std_logic_vector(4 downto 0) := "11111";
  constant st4: std_logic_vector(4 downto 0) := "10001";
  constant st5: std_logic_vector(4 downto 0) := "10110";
  constant st6: std_logic_vector(4 downto 0) := "01011";
  constant st7: std_logic_vector(4 downto 0) := "01111";
  constant st8: std_logic_vector(4 downto 0) := "00001";
  constant st9: std_logic_vector(4 downto 0) := "10000";
  constant st10: std_logic_vector(4 downto 0) := "11010";
  constant st11: std_logic_vector(4 downto 0) := "11000";
  constant st12: std_logic_vector(4 downto 0) := "01000";
  constant st13: std_logic_vector(4 downto 0) := "00100";
  constant st15: std_logic_vector(4 downto 0) := "01001";
  constant st14: std_logic_vector(4 downto 0) := "00110";
  constant st29: std_logic_vector(4 downto 0) := "11100";
  constant st31: std_logic_vector(4 downto 0) := "00011";
  constant st30: std_logic_vector(4 downto 0) := "10111";
  constant st17: std_logic_vector(4 downto 0) := "10011";
  constant st18: std_logic_vector(4 downto 0) := "10010";
  constant st19: std_logic_vector(4 downto 0) := "00111";
  constant st20: std_logic_vector(4 downto 0) := "01100";
  constant st21: std_logic_vector(4 downto 0) := "10101";
  constant st22: std_logic_vector(4 downto 0) := "10100";
  constant st23: std_logic_vector(4 downto 0) := "00000";
  constant st24: std_logic_vector(4 downto 0) := "01101";
  constant st25: std_logic_vector(4 downto 0) := "00101";
  constant st26: std_logic_vector(4 downto 0) := "11001";
  constant st27: std_logic_vector(4 downto 0) := "01010";
  constant st28: std_logic_vector(4 downto 0) := "01110";
  signal current_state, next_state: std_logic_vector(4 downto 0);
begin
  process(clock) begin
    if rising_edge(clock) then current_state <= next_state;
    end if;
  end process;
  process(input, current_state) begin
    next_state <= "-----"; output <= "---";
    case current_state is
      when st0 =>
        if std_match(input, "000000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st1; output <= "000";
        elsif std_match(input, "001000") then next_state <= st2; output <= "000";
        elsif std_match(input, "010000") then next_state <= st3; output <= "000";
        elsif std_match(input, "100000") then next_state <= st4; output <= "000";
        elsif std_match(input, "000101") then next_state <= st5; output <= "000";
        elsif std_match(input, "001001") then next_state <= st6; output <= "000";
        elsif std_match(input, "010001") then next_state <= st7; output <= "000";
        elsif std_match(input, "100001") then next_state <= st8; output <= "000";
        elsif std_match(input, "000110") then next_state <= st9; output <= "000";
        elsif std_match(input, "001010") then next_state <= st10; output <= "000";
        elsif std_match(input, "010010") then next_state <= st11; output <= "000";
        elsif std_match(input, "100010") then next_state <= st12; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st15; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st14; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st31; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st30; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st16 =>
        if std_match(input, "000000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st17; output <= "000";
        elsif std_match(input, "001000") then next_state <= st18; output <= "000";
        elsif std_match(input, "010000") then next_state <= st19; output <= "000";
        elsif std_match(input, "100000") then next_state <= st20; output <= "000";
        elsif std_match(input, "000101") then next_state <= st21; output <= "000";
        elsif std_match(input, "001001") then next_state <= st22; output <= "000";
        elsif std_match(input, "010001") then next_state <= st23; output <= "000";
        elsif std_match(input, "100001") then next_state <= st24; output <= "000";
        elsif std_match(input, "000110") then next_state <= st25; output <= "000";
        elsif std_match(input, "001010") then next_state <= st26; output <= "000";
        elsif std_match(input, "010010") then next_state <= st27; output <= "000";
        elsif std_match(input, "100010") then next_state <= st28; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st15; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st14; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st31; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st30; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st1 =>
        if std_match(input, "000000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st1; output <= "000";
        elsif std_match(input, "000010") then next_state <= st1; output <= "000";
        elsif std_match(input, "000011") then next_state <= st1; output <= "000";
        elsif std_match(input, "100011") then next_state <= st17; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st1; output <= "010";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st17 =>
        if std_match(input, "000000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st17; output <= "000";
        elsif std_match(input, "000010") then next_state <= st17; output <= "000";
        elsif std_match(input, "000011") then next_state <= st1; output <= "000";
        elsif std_match(input, "100011") then next_state <= st17; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st17; output <= "010";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st2 =>
        if std_match(input, "000000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st2; output <= "000";
        elsif std_match(input, "000010") then next_state <= st2; output <= "000";
        elsif std_match(input, "000011") then next_state <= st2; output <= "000";
        elsif std_match(input, "100011") then next_state <= st18; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st2; output <= "010";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st18 =>
        if std_match(input, "000000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st18; output <= "000";
        elsif std_match(input, "000010") then next_state <= st18; output <= "000";
        elsif std_match(input, "000011") then next_state <= st2; output <= "000";
        elsif std_match(input, "100011") then next_state <= st18; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st18; output <= "010";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st3 =>
        if std_match(input, "000000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st3; output <= "000";
        elsif std_match(input, "000010") then next_state <= st3; output <= "000";
        elsif std_match(input, "000011") then next_state <= st3; output <= "000";
        elsif std_match(input, "100011") then next_state <= st19; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st3; output <= "010";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st19 =>
        if std_match(input, "000000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st19; output <= "000";
        elsif std_match(input, "000010") then next_state <= st19; output <= "000";
        elsif std_match(input, "000011") then next_state <= st3; output <= "000";
        elsif std_match(input, "100011") then next_state <= st19; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st19; output <= "010";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st4 =>
        if std_match(input, "000000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st4; output <= "000";
        elsif std_match(input, "000010") then next_state <= st4; output <= "000";
        elsif std_match(input, "000011") then next_state <= st4; output <= "000";
        elsif std_match(input, "100011") then next_state <= st20; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st4; output <= "010";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st20 =>
        if std_match(input, "000000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st20; output <= "000";
        elsif std_match(input, "000010") then next_state <= st20; output <= "000";
        elsif std_match(input, "000011") then next_state <= st4; output <= "000";
        elsif std_match(input, "100011") then next_state <= st20; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st20; output <= "010";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st5 =>
        if std_match(input, "000001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000000") then next_state <= st5; output <= "000";
        elsif std_match(input, "000010") then next_state <= st5; output <= "000";
        elsif std_match(input, "000011") then next_state <= st5; output <= "000";
        elsif std_match(input, "100011") then next_state <= st21; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st5; output <= "010";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st21 =>
        if std_match(input, "000001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000000") then next_state <= st21; output <= "000";
        elsif std_match(input, "000010") then next_state <= st21; output <= "000";
        elsif std_match(input, "000011") then next_state <= st5; output <= "000";
        elsif std_match(input, "100011") then next_state <= st21; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st21; output <= "010";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st6 =>
        if std_match(input, "000001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000000") then next_state <= st6; output <= "000";
        elsif std_match(input, "000010") then next_state <= st6; output <= "000";
        elsif std_match(input, "000011") then next_state <= st6; output <= "000";
        elsif std_match(input, "100011") then next_state <= st22; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st6; output <= "010";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st22 =>
        if std_match(input, "000001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000000") then next_state <= st22; output <= "000";
        elsif std_match(input, "000010") then next_state <= st22; output <= "000";
        elsif std_match(input, "000011") then next_state <= st6; output <= "000";
        elsif std_match(input, "100011") then next_state <= st22; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st22; output <= "010";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st7 =>
        if std_match(input, "000001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000000") then next_state <= st7; output <= "000";
        elsif std_match(input, "000010") then next_state <= st7; output <= "000";
        elsif std_match(input, "000011") then next_state <= st7; output <= "000";
        elsif std_match(input, "100011") then next_state <= st23; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st7; output <= "010";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st23 =>
        if std_match(input, "000001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000000") then next_state <= st23; output <= "000";
        elsif std_match(input, "000010") then next_state <= st23; output <= "000";
        elsif std_match(input, "000011") then next_state <= st7; output <= "000";
        elsif std_match(input, "100011") then next_state <= st23; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st23; output <= "010";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st8 =>
        if std_match(input, "000001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000000") then next_state <= st8; output <= "000";
        elsif std_match(input, "000010") then next_state <= st8; output <= "000";
        elsif std_match(input, "000011") then next_state <= st8; output <= "000";
        elsif std_match(input, "100011") then next_state <= st24; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st8; output <= "010";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st24 =>
        if std_match(input, "000001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000000") then next_state <= st24; output <= "000";
        elsif std_match(input, "000010") then next_state <= st24; output <= "000";
        elsif std_match(input, "000011") then next_state <= st8; output <= "000";
        elsif std_match(input, "100011") then next_state <= st24; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st24; output <= "010";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st9 =>
        if std_match(input, "000010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st9; output <= "000";
        elsif std_match(input, "000000") then next_state <= st9; output <= "000";
        elsif std_match(input, "000011") then next_state <= st9; output <= "000";
        elsif std_match(input, "100011") then next_state <= st25; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st9; output <= "010";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st25 =>
        if std_match(input, "000010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st25; output <= "000";
        elsif std_match(input, "000000") then next_state <= st25; output <= "000";
        elsif std_match(input, "000011") then next_state <= st9; output <= "000";
        elsif std_match(input, "100011") then next_state <= st25; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st25; output <= "010";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st10 =>
        if std_match(input, "000010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st10; output <= "000";
        elsif std_match(input, "000000") then next_state <= st10; output <= "000";
        elsif std_match(input, "000011") then next_state <= st10; output <= "000";
        elsif std_match(input, "100011") then next_state <= st26; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st10; output <= "010";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st26 =>
        if std_match(input, "000010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st26; output <= "000";
        elsif std_match(input, "000000") then next_state <= st26; output <= "000";
        elsif std_match(input, "000011") then next_state <= st10; output <= "000";
        elsif std_match(input, "100011") then next_state <= st26; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st26; output <= "010";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st11 =>
        if std_match(input, "000010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st11; output <= "000";
        elsif std_match(input, "000000") then next_state <= st11; output <= "000";
        elsif std_match(input, "000011") then next_state <= st11; output <= "000";
        elsif std_match(input, "100011") then next_state <= st27; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st11; output <= "010";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st27 =>
        if std_match(input, "000010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st27; output <= "000";
        elsif std_match(input, "000000") then next_state <= st27; output <= "000";
        elsif std_match(input, "000011") then next_state <= st11; output <= "000";
        elsif std_match(input, "100011") then next_state <= st27; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st27; output <= "010";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st12 =>
        if std_match(input, "000010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000001") then next_state <= st12; output <= "000";
        elsif std_match(input, "000000") then next_state <= st12; output <= "000";
        elsif std_match(input, "000011") then next_state <= st12; output <= "000";
        elsif std_match(input, "100011") then next_state <= st28; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st12; output <= "010";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st28 =>
        if std_match(input, "000010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st28; output <= "000";
        elsif std_match(input, "000000") then next_state <= st28; output <= "000";
        elsif std_match(input, "000011") then next_state <= st12; output <= "000";
        elsif std_match(input, "100011") then next_state <= st28; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st28; output <= "010";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st13 =>
        if std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st13; output <= "100";
        elsif std_match(input, "000010") then next_state <= st13; output <= "100";
        elsif std_match(input, "000000") then next_state <= st13; output <= "100";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st29 =>
        if std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st29; output <= "100";
        elsif std_match(input, "000010") then next_state <= st29; output <= "100";
        elsif std_match(input, "000000") then next_state <= st29; output <= "100";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st15 =>
        if std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st15; output <= "000";
        elsif std_match(input, "000010") then next_state <= st15; output <= "000";
        elsif std_match(input, "000000") then next_state <= st15; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st15; output <= "011";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st31; output <= "011";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st31 =>
        if std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st31; output <= "000";
        elsif std_match(input, "000010") then next_state <= st31; output <= "000";
        elsif std_match(input, "000000") then next_state <= st31; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st15; output <= "011";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st0; output <= "000";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st31; output <= "011";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st16; output <= "000";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st14 =>
        if std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st14; output <= "000";
        elsif std_match(input, "000010") then next_state <= st14; output <= "000";
        elsif std_match(input, "000000") then next_state <= st14; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st0; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st0; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st0; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st0; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st0; output <= "000";
        elsif std_match(input, "000100") then next_state <= st0; output <= "000";
        elsif std_match(input, "001000") then next_state <= st0; output <= "000";
        elsif std_match(input, "010000") then next_state <= st0; output <= "000";
        elsif std_match(input, "100000") then next_state <= st0; output <= "000";
        elsif std_match(input, "000101") then next_state <= st0; output <= "000";
        elsif std_match(input, "001001") then next_state <= st0; output <= "000";
        elsif std_match(input, "010001") then next_state <= st0; output <= "000";
        elsif std_match(input, "100001") then next_state <= st0; output <= "000";
        elsif std_match(input, "000110") then next_state <= st0; output <= "000";
        elsif std_match(input, "001010") then next_state <= st0; output <= "000";
        elsif std_match(input, "010010") then next_state <= st0; output <= "000";
        elsif std_match(input, "100010") then next_state <= st0; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st14; output <= "001";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st30; output <= "001";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when st30 =>
        if std_match(input, "000011") then next_state <= st0; output <= "000";
        elsif std_match(input, "100011") then next_state <= st16; output <= "000";
        elsif std_match(input, "000001") then next_state <= st30; output <= "000";
        elsif std_match(input, "000010") then next_state <= st30; output <= "000";
        elsif std_match(input, "000000") then next_state <= st30; output <= "000";
        elsif std_match(input, "11--00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--100") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-00") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-100") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1100") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--101") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-01") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-101") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1101") then next_state <= st16; output <= "000";
        elsif std_match(input, "11--10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1-1-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "1--110") then next_state <= st16; output <= "000";
        elsif std_match(input, "-11-10") then next_state <= st16; output <= "000";
        elsif std_match(input, "-1-110") then next_state <= st16; output <= "000";
        elsif std_match(input, "--1110") then next_state <= st16; output <= "000";
        elsif std_match(input, "000100") then next_state <= st16; output <= "000";
        elsif std_match(input, "001000") then next_state <= st16; output <= "000";
        elsif std_match(input, "010000") then next_state <= st16; output <= "000";
        elsif std_match(input, "100000") then next_state <= st16; output <= "000";
        elsif std_match(input, "000101") then next_state <= st16; output <= "000";
        elsif std_match(input, "001001") then next_state <= st16; output <= "000";
        elsif std_match(input, "010001") then next_state <= st16; output <= "000";
        elsif std_match(input, "100001") then next_state <= st16; output <= "000";
        elsif std_match(input, "000110") then next_state <= st16; output <= "000";
        elsif std_match(input, "001010") then next_state <= st16; output <= "000";
        elsif std_match(input, "010010") then next_state <= st16; output <= "000";
        elsif std_match(input, "100010") then next_state <= st16; output <= "000";
        elsif std_match(input, "000111") then next_state <= st13; output <= "100";
        elsif std_match(input, "001011") then next_state <= st0; output <= "000";
        elsif std_match(input, "001111") then next_state <= st13; output <= "100";
        elsif std_match(input, "010011") then next_state <= st14; output <= "001";
        elsif std_match(input, "010111") then next_state <= st13; output <= "100";
        elsif std_match(input, "011011") then next_state <= st0; output <= "000";
        elsif std_match(input, "011111") then next_state <= st13; output <= "100";
        elsif std_match(input, "100111") then next_state <= st29; output <= "100";
        elsif std_match(input, "101011") then next_state <= st16; output <= "000";
        elsif std_match(input, "101111") then next_state <= st29; output <= "100";
        elsif std_match(input, "110011") then next_state <= st30; output <= "001";
        elsif std_match(input, "110111") then next_state <= st29; output <= "100";
        elsif std_match(input, "111011") then next_state <= st16; output <= "000";
        elsif std_match(input, "111111") then next_state <= st29; output <= "100";
        end if;
      when others => next_state <= "-----"; output <= "---";
    end case;
  end process;
end behaviour;
